`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:03:07 12/19/2021 
// Design Name: 
// Module Name:    C6_13_0 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module C6_13_0(
    input Load,
    input Count,
    input D0,
    input D1,
    input D2,
    input D3,
    input Clock,
    output Q0,
    output Q1,
    output Q2,
    output Q3,
    output CO
    );


endmodule
